`timescale 1ns / 1ps

module score(
    
    );
endmodule
